module tb();

reg clk,rst;
reg [7:0] x0_real,x1_real,x2_real,x3_real,x4_real,x5_real,x6_real,x7_real,x0_img,x1_img,x2_img,x3_img,x4_img,x5_img,x6_img,x7_img;
wire [7:0] y0_real,y1_real,y2_real,y3_real,y4_real,y5_real,y6_real,y7_real,y0_img, y1_img,y2_img,y3_img,y4_img,y5_img,y6_img,y7_img;

DIT_FFT dut(clk,rst,x0_real,x1_real,x2_real,x3_real,x4_real,x5_real,x6_real,x7_real,x0_img,x1_img,x2_img,x3_img,x4_img,x5_img,x6_img,x7_img,y0_real,y1_real,y2_real,y3_real,y4_real,y5_real,y6_real,y7_real,y0_img, y1_img,y2_img,y3_img,y4_img,y5_img,y6_img,y7_img);

initial begin
	clk=0;
	forever #5; clk=~clk;
end

initial begin
	x0_img=0;
	x1_img=0;
	x2_img=0;
	x3_img=0;
	x4_img=0;
	x5_img=0;
	x6_img=0;
	x7_img=0;
	x0_real=0;
	x1_real=0;
	x2_real=0;
	x3_real=0;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;
	#20
	x0_real=8'd1;
	x1_real=8'd1;
	x2_real=8'd1;
	x3_real=8'd1;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;	
	#200
	x7_real=8'd1;
	x6_real=8'd1;
	x5_real=8'd1;
	x4_real=8'd1;
	x3_real=0;
	x2_real=0;
	x1_real=0;
	x0_real=0;
	#200
	x0_real=0;
	x1_real=0;
	x2_real=0;
	x3_real=0;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;
	#20
	x7_real=8'd1;
	x6_real=8'd1;
	x5_real=8'd1;
	x4_real=8'd1;
	x0_real=8'd1;
	x1_real=8'd1;
	x2_real=8'd1;
	x3_real=8'd1;
	#200
	x0_real=0;
	x1_real=0;
	x2_real=0;
	x3_real=0;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;
	#20
	x7_real=8'd1;
	x6_real=8'd2;
	x5_real=8'd3;
	x4_real=8'd4;
	x0_real=8'd5;
	x1_real=8'd6;
	x2_real=8'd7;
	x3_real=8'd8;
	#400
	x0_real=0;
	x1_real=0;
	x2_real=0;
	x3_real=0;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;
	#20
	x7_real=8'd3;
	x6_real=8'd3;
	x5_real=8'd3;
	x4_real=8'd3;
	x0_real=8'd3;
	x1_real=8'd3;
	x2_real=8'd3;
	x3_real=8'd3;
	#400
	x0_real=0;
	x1_real=0;
	x2_real=0;
	x3_real=0;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;
	#20
	x7_real=8'd7;
	x6_real=8'd7;
	x5_real=8'd7;
	x4_real=8'd7;
	x0_real=8'd7;
	x1_real=8'd7;
	x2_real=8'd7;
	x3_real=8'd7;
	#400
	x0_real=0;
	x1_real=0;
	x2_real=0;
	x3_real=0;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;
	#20
	x7_real=8'd15;
	x6_real=8'd15;
	x5_real=8'd15;
	x4_real=8'd15;
	x0_real=8'd15;
	x1_real=8'd15;
	x2_real=8'd15;
	x3_real=8'd15;
	#600
	x0_real=0;
	x1_real=0;
	x2_real=0;
	x3_real=0;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;
	#20
	x7_real=8'd31;
	x6_real=8'd31;
	x5_real=8'd31;
	x4_real=8'd31;
	x0_real=8'd31;
	x1_real=8'd31;
	x2_real=8'd31;
	x3_real=8'd31;
	#800
	x0_real=0;
	x1_real=0;
	x2_real=0;
	x3_real=0;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;
	#20
	x7_real=8'd63;
	x6_real=8'd63;
	x5_real=8'd63;
	x4_real=8'd63;
	x0_real=8'd63;
	x1_real=8'd63;
	x2_real=8'd63;
	x3_real=8'd63;
	#800
	x0_real=0;
	x1_real=0;
	x2_real=0;
	x3_real=0;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;
	#20
	x7_real=8'd127;
	x6_real=8'd127;
	x5_real=8'd127;
	x4_real=8'd127;
	x0_real=8'd127;
	x1_real=8'd127;
	x2_real=8'd127;
	x3_real=8'd127;
	#1000
	x0_real=0;
	x1_real=0;
	x2_real=0;
	x3_real=0;
	x4_real=0;
	x5_real=0;
	x6_real=0;
	x7_real=0;
	#20
	x7_real=8'd1;
	x6_real=8'd1;
	x5_real=8'd1;
	x4_real=8'd1;
	x0_real=8'd1;
	x1_real=8'd1;
	x2_real=8'd1;
	x3_real=8'd1;
end

endmodule
